-- this circuit converts a 6-bit binary number to a 2-digit BCD representation --
-- entity name: g01_binary_to_BCD 
--
-- Copyright (C) 2014 Alex Carruthers, Dan Grencorn 
-- Version 1.0
-- Author: Alex Carruthers, Dan Greencorn; michael.carruthers@mail.mcgill.ca, dan.greencorn@mail.mcgill.ca 
-- Date: February 13, 2014

library ieee; 
-- allows use of the std_logic_vector type
use ieee.std_logic_1164.all;
use ieee.numeric_std.all; -- allows use of the unsigned type

library lpm; -- allows use of the Altera library modules 
use lpm.lpm_components.all;

entity g01_binary_to_BCD is
	port ( clock : in std_logic; -- to clock the lpm_rom register
		bin : in unsigned(5 downto 0);
		BCD : out std_logic_vector(7 downto 0)
	);
end g01_binary_to_BCD;

architecture converter of g01_binary_to_BCD is

begin
	bcd_table : lpm_rom
		GENERIC MAP(
			lpm_widthad => 6,
			lpm_numwords => 64,
			lpm_outdata => "UNREGISTERED",
			lpm_address_control => "REGISTERED",
			lpm_file => "g01_binary_to_BCD.mif",
			lpm_width => 8
		)
		PORT MAP (clock => clock, address => bin, q => BCD);
end converter;